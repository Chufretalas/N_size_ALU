PACKAGE my_types IS
    TYPE T_Operations IS (OP_AND, OP_OR, OP_Adder, OP_Less);
END PACKAGE;